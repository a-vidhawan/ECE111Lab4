// 2to1 Multiplexor behavioral code
module mux_2x1(
  input in0, in1, 
  input sel, 
  output logic out
); 

// fill in the guts
//  pseudocode: out =sel? in1 : in0;
endmodule
 

